entity lab4 is
	port(clock : in bit)